// Copyright 2022 Sabana Technologies, Inc
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module sabana (
  input  logic clock,
  input  logic reset,
  input  logic start,
  output logic finish,
  input  logic [32-1:0] a_in,
  input  logic [32-1:0] b_in,
  input  logic [32-1:0] c_in,
  output logic [32-1:0] y_out,
  output logic y_valid
);

  logic is_finish;
  always_ff @(posedge clock)
    if (reset)
      is_finish <= 1'b0;
    else
      is_finish <= start;

  toplevel toplevel_i (
    .clock(clock),
    .rst(reset),
    .a(a_in),
    .b(b_in),
    .c(c_in),
    .y(y_out)
  );

  assign y_valid = is_finish;
  assign finish = is_finish;

endmodule
